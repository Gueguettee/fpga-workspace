

architecture arch of task5 is
    