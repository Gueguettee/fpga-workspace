library ieee;
use ieee.std_logic_1164.all;

package my_pkg is 
	constant DATA_BUS_WIDTH_c : integer := 32;

end my_pkg;